
-------------------------------------------------------
--! @file
--! @brief PONG Hauptentity 
-------------------------------------------------------
entity PONG is
    port(
        clk: in bit
    );
end entity;


architecture PONG_ARC of PONG is


begin


end architecture;
