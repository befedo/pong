library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity VGA_RAM is    
	generic(
        --! Horizontale groesse des Rams.
       H_WIDTH:natural:=8;
        --! Vertikale groesse des Rams.
       V_WIDTH:natural:=8;
        --! Breite eines Speicherbereichs.
       WORD_WIDTH:natural:=3
    );
    port(
        --! Adresseingang fr die Horizontale.
        H_ADR: in std_logic_vector(H_WIDTH-1 downto 0);
        --! Adresseingang fr die Vertikale.
        V_ADR: in std_logic_vector(V_WIDTH-1 downto 0);
        --! Eingangsleitung zum Parallelen schreiben.
        DIN: in std_logic_vector(WORD_WIDTH-1 downto 0);
        --! Alle Operationen werden mit denn Takt synchronisiert.
        CLK: in std_logic;
        --! Wenn das signal High ist wird das aktuelle Signal am DIN gespeichert. EN muss auch HIGH sein damit ein Effekt auftritt.
        WE: in std_logic;
        --! Wenn das signal High ist wird der Speicherbaustein aktiv.
        EN: in std_logic;
        --! Datenausgangsleitung zum Parallelen lesen.
        DOUT: out std_logic_vector(WORD_WIDTH-1 downto 0)
    );
end entity VGA_RAM;

architecture VGA_RAM_ARC of VGA_RAM is
type MEM is array (0 to 2**(H_WIDTH+V_WIDTH)-1) of std_logic_vector(WORD_WIDTH-1 downto 0);
signal MEM_MAIN: MEM:=(	"100","010","001","010","111","110","101","101","101","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","111","010","100","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						"111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010","111","110","001","010",
						
						others=>"000");
signal ADR: std_logic_vector(H_WIDTH+V_WIDTH-1 downto 0);
begin


    process(CLK,EN)
    begin
        if(EN= '1' ) then
            if (CLK'Event and CLK = '1') then
                                ADR(V_WIDTH-1 downto 0)<=V_ADR;
                                ADR(H_WIDTH+V_WIDTH-1 downto V_WIDTH)<=H_ADR;
                if(WE = '1' ) then
                    MEM_MAIN(to_integer(unsigned(ADR)))<=DIN;
                end if;
            end if;
        end if;
    end process;
    
    DOUT<=MEM_MAIN(to_integer(unsigned(ADR)));

end architecture VGA_RAM_ARC;